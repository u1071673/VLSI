
module i2c (
	input wire clk,
	input wire rst,
	output reg sda,
	output reg scl
	);
endmodule
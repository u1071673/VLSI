
module seven_segment_controller (
	input clk,    // Clock
	input rst,
	input hundreds,
	input tens,
	input ones,
	output a,
	output b,
	output c,
	output d,
	output e,
	output f,
	output g
);

endmodule

module pad_out_buffered(
	input out,
	output pad
);

INVX1 inv0 (.A(out), .Z(out_pre));
INVX4 inv1 (.A(out_pre), .Z(out_pre1));
INVX16 inv2 (.A(out_pre1), .Z(out_pre2));
INVX32 inv3 (.A(out_pre2), .Z(out_buf));
pad_out pad_out0(.pad(pad), .DataOut(out_buf));
endmodule // pad_out_buffered
